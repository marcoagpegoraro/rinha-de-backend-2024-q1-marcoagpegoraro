module dtos

pub struct TransacaoResponseDto {
pub:
	limite 	i64
	saldo 	i64
}
