module main

fn main(){
	print("Hello, world")
}